//Simulation File

`timescale 1ns / 1ps

interface full_adder_if;
    
    logic A;
    logic B;
    logic Cin;
    logic SUM;
    logic CARRY;

endinterface