//Simulation file

`timescale 1ns / 1ps

interface half_adder_if;
    
    logic A;
    logic B;
    logic SUM;
    logic CARRY;
    
endinterface
